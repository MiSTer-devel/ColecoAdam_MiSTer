`timescale 1ns / 1ps

module sdpramv #(
    parameter widthad_a = 10,
    parameter width_a = 8,
    parameter init_file= ""
) (
    input   wire                clock,
    input   wire                wren_a,
    input   wire    [widthad_a-1:0]  address_a,
    input   wire    [width_a-1:0]  data_a,
    output  reg     [width_a-1:0]  q_a,
    input   wire                wren_b,
    input   wire    [widthad_a-1:0]  address_b,
    input   wire    [width_a-1:0]  data_b,
    output  reg     [width_a-1:0]  q_b,

    input wire cs,
    input wire enable
);

    initial begin
        $display("Loading rom.");
        $display(init_file);
        if (init_file>0)
                $readmemh(init_file, mem);
    end


// Shared memory
reg [width_a-1:0] mem [(2**widthad_a)-1:0];

always @(posedge clock) begin
    q_a      <= mem[address_a];
    q_b      <= mem[address_b];
    if(wren_a) begin
//$display("writing %x %x",address,data);
        q_a      <= data_a;
        mem[address_a] <= data_a;
    end
    if(wren_b) begin
//$display("writing %x %x",address,data);
        q_b      <= data_b;
        mem[address_b] <= data_b;
    end
end


endmodule
